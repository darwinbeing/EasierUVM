covergroup m_cov;
  option.per_instance = 1;
  cp_data: coverpoint m_item.data;
endgroup
