package common_pkg;
endpackage
