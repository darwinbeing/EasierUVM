function void refmodel::write_refmodel_0(mytrans t);                                                  

endfunction                                                                                      
