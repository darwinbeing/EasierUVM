typedef struct packed {
  bit cmd;
  byte addr;
  byte data;
} bus_tx_s;
