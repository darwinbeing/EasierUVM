package common_env_pkg;
endpackage
