  extern function new(string name, uvm_component parent);
  extern function void write(input bus_tx t);
  extern function void build_phase(uvm_phase phase);
