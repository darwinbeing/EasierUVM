covergroup m_cov;
  option.per_instance = 1;
  coverpoint m_item.data;
endgroup: m_cov
