extern task          run_phase(uvm_phase phase);

extern function void write(bus_tx_s req_s);
