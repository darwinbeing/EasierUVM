module dut;

endmodule
